-- altera vhdl_input_version vhdl_2008

-- Lucas Ritzdorf
-- 04/30/2024
-- EELE 468

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-- HPS interface for convolution processor
entity convolutionProcessor is
    port (
        clk                      : in  std_logic;  -- system clock
        reset                    : in  std_logic;  -- system reset, active high

        -- Avalon streaming interface (audio sink)
        avalon_st_sink_valid     : in  std_logic;
        avalon_st_sink_data      : in  std_logic_vector(23 downto 0);
        avalon_st_sink_channel   : in  std_logic_vector(0 downto 0);
        -- Avalon streaming interface (audio source)
        avalon_st_source_valid   : out std_logic;
        avalon_st_source_data    : out std_logic_vector(23 downto 0);
        avalon_st_source_channel : out std_logic_vector(0 downto 0);

        -- Avalon memory-mapped interface (control registers)
        avalon_mm_address        : in  std_logic_vector(1 downto 0);
        avalon_mm_read           : in  std_logic;
        avalon_mm_readdata       : out std_logic_vector(31 downto 0);
        avalon_mm_write          : in  std_logic;
        avalon_mm_writedata      : in  std_logic_vector(31 downto 0);

        -- Real-time control signals
        rt_record                : in  std_logic;
        rt_recording             : out std_logic;
        rt_enabled               : out std_logic
    );
end entity;


architecture convolutionProcessor_Arch of convolutionProcessor is

    -- Actual convolution component, generated by MATLAB HDL Coder
    component convolutionPlayback is
        port (
            clk         : in    std_logic;
            reset       : in    std_logic;
            clk_enable  : in    std_logic;
            audioIn     : in    std_logic_vector(23 downto 0);
            modeControl : in    std_logic;
            wetDryMix   : in    std_logic_vector(15 downto 0);
            volume      : in    std_logic_vector(15 downto 0);
            enable      : in    std_logic;
            ce_out      : out   std_logic;
            audioOut    : out   std_logic_vector(23 downto 0);
            recording   : out   std_logic
        );
    end component;

    -- Avalon streaming to left/right-clocked interface converter
    component ast2lr is
        port (
            clk                 : in  std_logic;
            avalon_sink_data    : in  std_logic_vector(23 downto 0);
            avalon_sink_channel : in  std_logic;
            avalon_sink_valid   : in  std_logic;
            data_left           : out std_logic_vector(23 downto 0);
            data_right          : out std_logic_vector(23 downto 0)
        );
    end component ast2lr;

    -- Left/right-clocked to Avalon streaming interface converter
    component lr2ast is
        port (
            clk                   : in  std_logic;
            avalon_sink_channel   : in  std_logic;
            avalon_sink_valid     : in  std_logic;
            data_left             : in  std_logic_vector(23 downto 0);
            data_right            : in  std_logic_vector(23 downto 0);
            avalon_source_data    : out std_logic_vector(23 downto 0);
            avalon_source_channel : out std_logic;
            avalon_source_valid   : out std_logic
        );
    end component lr2ast;

    -- Internal audio data signals
    signal
        left_sink_data, right_sink_data,
        left_source_data, right_source_data
        : std_logic_vector(23 downto 0);

    -- Avalon-mapped control registers
    -- NOTE: These apply to both channels (i.e. mono control), though stereo
    --     control is achievable by duplicating the registers and connecting
    --     them to the appropriate component instances.
    signal wetDryMix : std_logic_vector(15 downto 0);  -- UQ0.16
    signal volume    : std_logic_vector(15 downto 0);  -- UQ0.16
    signal enable    : std_logic;
    signal left_recording, right_recording : std_logic;

begin

    u_ast2lr : component ast2lr
        port map (
            clk                 => clk,
            avalon_sink_data    => avalon_st_sink_data,
            avalon_sink_channel => avalon_st_sink_channel(0),
            avalon_sink_valid   => avalon_st_sink_valid,
            data_left           => left_sink_data,
            data_right          => right_sink_data
        );
    u_lr2ast : component lr2ast
        port map (
            clk                   => clk,
            avalon_sink_channel   => avalon_st_sink_channel(0),
            avalon_sink_valid     => avalon_st_sink_valid,
            data_left             => left_source_data,
            data_right            => right_source_data,
            avalon_source_data    => avalon_st_source_data,
            avalon_source_channel => avalon_st_source_channel(0),
            avalon_source_valid   => avalon_st_source_valid
        );

    -- One filter system for each channel
    left_filter : component convolutionPlayback
        port map (
            clk         => clk,
            reset       => reset,
            clk_enable  => '1',
            audioIn     => left_sink_data,
            modeControl => rt_record,
            wetDryMix   => wetDryMix,
            volume      => volume,
            enable      => enable,
            ce_out      => open,
            audioOut    => left_source_data,
            recording   => left_recording
        );
    right_filter : component convolutionPlayback
        port map (
            clk         => clk,
            reset       => reset,
            clk_enable  => '1',
            audioIn     => right_sink_data,
            modeControl => rt_record,
            wetDryMix   => wetDryMix,
            volume      => volume,
            enable      => enable,
            ce_out      => open,
            audioOut    => right_source_data,
            recording   => right_recording
        );

    -- Manage reading from mapped registers
    avalon_register_read : process (clk) is
    begin
        if rising_edge(clk) and (?? avalon_mm_read) then
            case avalon_mm_address is
                when "00" => avalon_mm_readdata <= std_logic_vector(resize(unsigned(wetDryMix), avalon_mm_readdata'length));
                when "01" => avalon_mm_readdata <= std_logic_vector(resize(unsigned(volume   ), avalon_mm_readdata'length));
                when "10" => avalon_mm_readdata <= std_logic_vector(to_unsigned(0, avalon_mm_readdata'length-1)) & enable;
                when others => null;
            end case;
        end if;
    end process;

    -- Manage writing to mapped registers
    avalon_register_write : process (clk, reset) is
    begin
        if reset then
            wetDryMix <= "1111111111111111";  -- All "wet", no "dry" signal
            volume    <= "1000000000000000";  -- One-half
            enable    <= '1';
        elsif rising_edge(clk) and (?? avalon_mm_write) then
            case avalon_mm_address is
                when "00" => wetDryMix <= std_logic_vector(resize(unsigned(avalon_mm_writedata), wetDryMix'length));
                when "01" => volume    <= std_logic_vector(resize(unsigned(avalon_mm_writedata), volume'length));
                when "10" =>
                    -- This should be a one-liner, but Quartus doesn't like the unary "or" operator
                    if avalon_mm_writedata /= std_logic_vector(to_unsigned(0, avalon_mm_readdata'length)) then
                        enable <= '1';
                    else
                        enable <= '0';
                    end if;
                when others => null;
            end case;
        end if;
    end process;

    -- Assign real-time output signals
    rt_recording <= left_recording or right_recording;
    rt_enabled <= enable;

end architecture;
